/*********************************************************
 MODULE:        Sub Level SDRAM Refresh Acknowledge

 FILE NAME:    ref_ack.v
 VERSION:    1.0
 DATE:        April 28th, 2002
 AUTHOR:        Hossein Amidi
 COMPANY:    
 CODE TYPE:    Register Transfer Level

 DESCRIPTION:    This module is the sub level RTL code of SDRAM Controller ASIC verilog
 code. It is the Refresh Acknowledge block.


 Hossein Amidi
 (C) April 2002

*********************************************************/

// DEFINES
`timescale 1ns / 10ps

module ref_ack(// Input
                    reset,
                    clk0,
                    do_refresh,
                    do_reada,
                    do_writea,
                    do_preacharge,
                    do_load_mod,
                    ref_req,
                    // Output
                    cmack,
                    ref_ack
                    );

// Parameter
`include        "parameter.v"

// Input
input reset;
input clk0;
input do_refresh;
input do_reada;
input do_writea;
input do_preacharge;
input do_load_mod;
input ref_req;

// Output
output cmack;
output ref_ack;

// Internal wire and reg signals
wire reset;
wire clk0;
wire do_refresh;
wire do_reada;
wire do_writea;
wire do_preacharge;
wire do_load_mod;
wire ref_req;

reg    cmack;
reg   ref_ack;

// Assignment

// This always block generates the command acknowledge, cmack, signal.
// It also generates the acknowledge signal, ref_ack, that acknowledges
// a refresh request that was generated by the internal refresh timer circuit.
always @(posedge reset or posedge clk0) 
begin

        if (reset == 1'b1) 
        begin
                cmack    <= 0;
                ref_ack  <= 0;
        end
        
        else
        begin
                if (do_refresh == 1 & ref_req == 1)                   // Internal refresh timer refresh request
                        ref_ack <= 1;
                else if ((do_refresh == 1) | (do_reada == 1) | (do_writea == 1) | (do_preacharge == 1)   // externa  commands
                         | (do_load_mod))
                        cmack <= 1;
                else
                begin
                        ref_ack <= 0;
                        cmack   <= 0;
                end
        end
end 


endmodule
